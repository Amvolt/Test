module delay(DelayTime);
